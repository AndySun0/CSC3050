`timescale 1ns / 10ps
`include "./ALU.v"
`include "./Signal.v"
`include "./stages.v"


module PC_checker(CLK, NEW_PC, BRC_PC, PC_BRCH_INTO, JUMP_TO_PC, JUMPSIGN, PC_write, PC);
    input CLK, PC_BRCH_INTO, PC_write, JUMPSIGN;
    input [31:0] NEW_PC, BRC_PC, JUMP_TO_PC;
    output reg [31:0] PC;

    initial
    PC = 32'b0;
    
    always @(posedge CLK) begin
        if (PC_write) begin
            if (PC_BRCH_INTO) begin
                PC <= BRC_PC;
            end else if (JUMPSIGN) begin
                PC <= JUMP_TO_PC;
            end else begin
                PC <= NEW_PC;
            end
        end else if (~PC_write) begin
            PC <= NEW_PC - 4;
        end
    end
    endmodule


module instruction_memory (CLK , PC , ENABLE , NEW_PC , INSTRUCTION);
    input CLK , ENABLE;
    input[31:0] PC;
    output reg[31:0] NEW_PC , INSTRUCTION;

    reg[31:0] RAM[0:512-1];
    initial begin
    $readmemb("CPU_instruction.bin", RAM);
    end

    always @(PC) begin               // when instruction_pc changes to a new value, the INSTRUCTION memory can fetch the target instrucion
        if(ENABLE == 1) begin
            INSTRUCTION <= RAM[PC/4];    // if ENABLE == 1 it means the INSTRUCTION memory can work at this time
            NEW_PC <= PC + 4;            // at the same time add PC and 4 to get the potential next INSTRUCTION palce
        end
        
    end
endmodule

module enable_checker (INSTRUCTION , ENABLE);
    input[31:0] INSTRUCTION;
    output reg ENABLE;
    initial begin
        ENABLE = 1;
    end
    always @(INSTRUCTION) begin
        // if(INSTRUCTION == 32'b11111111111111111111111111111111) begin
        //     ENABLE <= 1'b0;
        // end
        // else begin
        //     ENABLE <= 1'b1;
        case (INSTRUCTION) 
            32'b1111_1111_1111_1111_1111_1111_1111_1111:
            ENABLE <= 1'b0;
            default:
            ENABLE <= 1'b1;
        endcase
        end
    
endmodule

// module IF_ID_buffer(INSTRUCTION , NEW_PC , IF_flush , IF_ID_write , CLK , ENABLE , next_PC , instruction_F);
//     input[31:0] INSTRUCTION , NEW_PC;
//     input IF_flush , IF_ID_write , CLK , ENABLE;
//     output reg[31:0] next_PC , instruction_F;

//     always @(posedge CLK) begin
//         if (ENABLE == 1) begin
//             if(IF_flush == 1) begin
//                 next_PC <= NEW_PC;
//                 instruction_F <= 0;
//             end
//             else if(IF_ID_write == 1) begin
//                 next_PC <= NEW_PC;
//                 instruction_F <= INSTRUCTION;
//             end
//             else if(IF_ID_write == 0) begin
//                 next_PC <= next_PC;
//                 instruction_F <= instruction_F;
//             end
//         end
//     end
// endmodule

module decode (instruction_F , opcode , rs , rt , rd , imme , funct , shamt , target);
    input[31:0] instruction_F;
    output reg[5:0] opcode;
    output reg[4:0] rs , rt , rd , shamt;
    output reg[15:0] imme;
    output reg[5:0] funct;
    output reg[25:0] target;

    always @(instruction_F) begin
        opcode <= instruction_F[31:26];
        rs <= instruction_F[25:21];
        rt <= instruction_F[20:16];
        rd <= instruction_F[15:11];
        shamt <= instruction_F[10:6];
        funct <= instruction_F[5:0];
        imme <= instruction_F[15:0];
        target <= instruction_F[25:0];
    end
endmodule


module Register (CLK , next_PC , write_back_data , write_registerW , RegwriteW , opcode , rs , rt , imme ,
                 target , read_data1 , read_data2 , BRC_PC , JUMP_TO_PC , zero_flag);
    input CLK , RegwriteW;
    input[31:0] next_PC , write_back_data;
    input[5:0] opcode;
    input[4:0] write_registerW , rs , rt;
    input[15:0] imme;
    input[25:0] target;
    output reg[31:0] read_data1 , read_data2;
    output reg[31:0] BRC_PC , JUMP_TO_PC;
    output reg zero_flag;
    reg[31:0] ext_imme;
    reg[31:0] Reg[0:31];

    integer i;
    initial begin
        for (i=0; i < 32; i = i + 1) begin
            Reg[i] = 32'b0;
        end
    end

    always @(posedge CLK) begin  //write in data in the first half clock write_registerW
        if(RegwriteW == 1)begin
            Reg[write_registerW] <= write_back_data;
        end
    end

    always @(negedge CLK) begin  //read data out in the second half clock
        read_data1 <= Reg[rs];
        read_data2 <= Reg[rt];
    end

    // always @(read_data2 , read_data1) begin
    //     case(opcode)
    //     6'b000100: begin          //beq function
    //         if(read_data1 == read_data2) begin
    //             zero_flag <= 1;
    //         end 
    //         else begin
    //             zero_flag <= 0;
    //         end
    //     end
    //     6'b000101: begin          //bne function
    //         if(read_data1 == read_data2) begin
    //             zero_flag <= 0;
    //         end 
    //         else begin
    //             zero_flag <= 1;
    //         end
    //     end
    //     default: zero_flag <= 0;
    //     endcase
    // end
    always @* begin
        case (opcode)
            6'b000100: zero_flag <= (read_data1 == read_data2);
            6'b000101: zero_flag <= (read_data1 != read_data2);
            default: zero_flag <= 0;
        endcase
    end

    // always @(imme) begin        //extend the imme number accorfing to the INSTRUCTION requirment
    //     ext_imme <= $signed(imme);
    // end

    // always @(ext_imme) begin    //calculate the branch PC after the extimme is ready
    //     BRC_PC = next_PC + ext_imme * 4;
    // end

    // always @(read_data1 , target , opcode) begin
    //     case (opcode)
    //         6'b000000: begin
    //             JUMP_TO_PC <= read_data1;
    //         end
    //         6'b000010: begin
    //             JUMP_TO_PC <= target * 4;
    //         end
    //         6'b000011: begin
    //             JUMP_TO_PC <= target * 4;
    //         end
    //         default: JUMP_TO_PC <= 0;
    //     endcase
    // end
    always @* begin
        ext_imme = $signed(imme);
    end

    always @* begin
        BRC_PC = next_PC + ext_imme * 4;
    end

    always @* begin
        case (opcode)
            6'b000000: JUMP_TO_PC <= read_data1;
            6'b000010, 6'b000011: JUMP_TO_PC <= target * 4;
            default: JUMP_TO_PC <= 0;
        endcase
    end

endmodule

// module hazard_unit (rs , rt , rt_E , MemreadE , MemwriteE , PC_write , IF_ID_write , ID_EX_flush);
//     input[4:0] rs , rt , rt_E;
//     input MemreadE , MemwriteE;
//     output reg PC_write , IF_ID_write , ID_EX_flush;
//     initial begin
//         PC_write = 1;
//         IF_ID_write = 1;
//     end
//     always @(rs , rt , rt_E , MemreadE , MemwriteE) begin
//         if((MemreadE & (rt_E == rt)) || (MemreadE & (rt_E == rs))) begin         //lw instructions will cause hazard
//             PC_write <= 0;
//             IF_ID_write <= 0;
//             ID_EX_flush <= 0;
//         end
//         else if((MemwriteE & (rt_E == rt)) || (MemwriteE & (rt_E == rs))) begin
//             PC_write <= 0;
//             IF_ID_write <= 0;
//             ID_EX_flush <= 0;
//         end
//         else begin
//             PC_write <= 1;
//             IF_ID_write <= 1;
//             ID_EX_flush <= 1;
//         end
//     end
// endmodule
module hazard_unit (rs , rt , rt_E , MemreadE , MemwriteE , PC_write , IF_ID_write , ID_EX_flush);
    input[4:0] rs , rt , rt_E;
    input MemreadE , MemwriteE;
    output reg PC_write , IF_ID_write , ID_EX_flush;
    always @* begin
        if((MemreadE && (rt_E == rt || rt_E == rs)) ||
        (MemwriteE && (rt_E == rt || rt_E == rs))) begin
            PC_write = 0;
            IF_ID_write = 0;
            ID_EX_flush = 0;
        end
        else begin
            PC_write = 1;
            IF_ID_write = 1;
            ID_EX_flush = 1;
        end
    end

    initial begin
        PC_write = 1;
        IF_ID_write = 1;
        ID_EX_flush = 0;
    end
endmodule

// module ID_EX_buffer (
//     input CLK,
//     input [31:0] read_data1,
//     input [31:0] read_data2,
//     input [5:0] opcode,
//     input [4:0] rs,
//     input [4:0] rt,
//     input [4:0] rd,
//     input [15:0] imme,
//     input [25:0] target,
//     input [4:0] shamt,
//     input [5:0] funct,
//     input RegDstD,
//     input MemreadD,
//     input MemtoRegD,
//     input [2:0] ALUopD,
//     input MemwriteD,
//     input ALUSrcD,
//     input RegwriteD,
//     input sign_extD,
//     output reg [31:0] read_data_E1,
//     output reg [31:0] read_data_E2,
//     output reg [5:0] opcode_E,
//     output reg [4:0] rs_E,
//     output reg [4:0] rt_E,
//     output reg [4:0] rd_E,
//     output reg [15:0] imme_E,
//     output reg [25:0] target_E,
//     output reg [4:0] shamt_E,
//     output reg [5:0] funct_E,
//     output reg RegDstE,
//     output reg MemreadE,
//     output reg MemtoRegE,
//     output [2:0] ALUopE,
//     output reg MemwriteE,
//     output reg ALUSrcE,
//     output reg RegwriteE,
//     output reg sign_extE,
//     output reg [31:0] next_PC_E
//     );
    
    // always @(posedge CLK) begin
    //     read_data_E1 <= read_data1;
    //     read_data_E2 <= read_data2;
    //     imme_E <= imme;
    //     opcode_E <= opcode;
    //     shamt_E <= shamt;
    //     funct_E <= funct;
    //     rs_E <= rs;
    //     rt_E <= rt;
    //     rd_E <= rd;
    //     RegDstE <= RegDstD;
    //     MemreadE <= MemreadD;
    //     MemtoRegE <= MemtoRegD;
    //     ALUopE <= ALUopD;
    //     MemwriteE <= MemwriteD;
    //     ALUSrcE <= ALUSrcD;
    //     RegwriteE <= RegwriteD;
    //     sign_extE <= sign_extD;
    //     target_E <= target;
    //     next_PC_E <= next_PC;
    // end


module Write_register_checker (opcode_E , rt_E , rd_E , RegDstE , write_register);
    input[4:0] rt_E , rd_E;
    input[5:0] opcode_E;
    input RegDstE;
    output reg[4:0]write_register;
    always @(opcode_E , rt_E , rd_E , RegDstE) begin
        if(opcode_E == 6'b000011) 
            write_register = 5'b11111;
        // end
        // else begin
        //     if(RegDstE == 0) write_register = rt_E;
        //     else if (RegDstE == 1) write_register = rd_E;
        else if (RegDstE == 0)
            write_register = rt_E;
        else if (RegDstE == 1)
            write_register = rd_E;
        
        end
endmodule

module forwarding_unit (CLK , rs_E , rt_E , write_registerM , write_registerW , RegwriteM , RegwriteW , rs_source , rt_source);
    input[4:0] rs_E , rt_E , write_registerM , write_registerW;
    input RegwriteM , RegwriteW , CLK;
    output reg[1:0] rs_source , rt_source;
    always @(rs_E , rt_E , write_registerM , write_registerW , RegwriteM , RegwriteW , posedge CLK) begin
        if(RegwriteM == 1 && write_registerM != 0 && write_registerM == rs_E)begin
            rs_source <= 2'b10;
        end
        else if(RegwriteW == 1 && write_registerW != 0 && write_registerW == rs_E) begin
            rs_source <= 2'b01;
        end
        else begin
            rs_source <= 2'b00;
        end
        if(RegwriteM == 1 && write_registerM != 0 && write_registerM == rt_E)begin
            rt_source <= 2'b10;
        end
        else if(RegwriteW == 1 && write_registerW != 0 && write_registerW == rt_E) begin
            rt_source <= 2'b01;
        end
        else begin
            rt_source <= 2'b00;
        end
    end
    // always @(posedge CLK) begin
    //     if (RegwriteM == 1 && write_registerM != 0 && write_registerM == rs_E) begin
    //         rs_source <= 2'b10;
    //     end else if (RegwriteW == 1 && write_registerW != 0 && write_registerW == rs_E) begin
    //         rs_source <= 2'b01;
    //     end else begin
    //         rs_source <= 2'b00;
    //     end
        
    //     if (RegwriteM == 1 && write_registerM != 0 && write_registerM == rt_E) begin
    //         rt_source <= 2'b10;
    //     end else if (RegwriteW == 1 && write_registerW != 0 && write_registerW == rt_E) begin
    //         rt_source <= 2'b01;
    //     end else begin
    //         rt_source <= 2'b00;
    //     end
    // end

endmodule

module Check_write_back_data (MemtoRegW , ALU_resultW , MemdataW , write_back_data);
    input MemtoRegW;
    input[31:0] ALU_resultW , MemdataW;
    output reg[31:0] write_back_data;

    always @(MemtoRegW , ALU_resultW , MemdataW) begin
        if(MemtoRegW == 0) begin
            write_back_data <= ALU_resultW;
        end
        else if(MemtoRegW == 1) begin
            write_back_data <= MemdataW;
        end
    end
endmodule

module MainMemory (ALU_resultM , write_dataM , MemreadM , MemwriteM , Memdata);
    input[31:0] ALU_resultM , write_dataM;
    input MemreadM , MemwriteM;
    output reg[31:0] Memdata;

    reg [31:0] DATA_RAM [0:512-1];

    reg [16383:0] ram_init;
    integer i;
    initial begin
        ram_init = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
        for (i=0; i < 512; i = i + 1) begin
            DATA_RAM[512-1-i] = ram_init[i*32+:32];
        end
    end

    always @(MemreadM , MemwriteM , write_dataM , ALU_resultM) begin
        if(MemreadM == 1)begin
            Memdata <= DATA_RAM[ALU_resultM/4];
        end
        else if(MemwriteM == 1)begin
            DATA_RAM[ALU_resultM/4] <= write_dataM;
            //$display("write %b in %b", write_dataM, ALU_resultM/4);
            Memdata <= 0;
        end
        else Memdata <= 0;
    end
endmodule

module CPU(
    input wire CLK
    );
    // reg CLK;
    reg[31:0] pc;
    // initial CLK = 1'b0;
    // always #5 CLK = ~CLK;
    wire ENABLE;
    wire PC_write;
    wire[31:0] PC;
    wire[31:0] BRC_PC;
    wire[31:0] NEW_PC;
    wire[31:0] INSTRUCTION;
    wire IF_flush;
    wire IF_ID_write = 1'b1;
    wire[31:0] next_PC;
    wire[31:0] instruction_F;
    wire[5:0] opcode;
    wire[4:0] rs , rt , rd , shamt;
    wire[15:0] imme;
    wire[5:0] funct;
    wire[25:0] target;
    wire ID_EX_flush , zero_flag;
    wire RegDst , Branch , Memread , MemtoReg , ALUop , Memwrite , ALUSrc , Regwrite , sign_ext , PC_BRCH_INTO , JUMPSIGN;
    wire[31:0] write_back_data;
    wire[31:0] read_data1 , read_data2;
    wire[31:0] JUMP_TO_PC;
    wire[15:0] imme_E;
    wire[31:0] read_data_E1 , read_data_E2 , next_PC_E;
    wire[5:0] opcode_E , funct_E;
    wire[4:0] rs_E , rt_E , rd_E , shamt_E;
    wire RegDstE , MemreadE , MemtoRegE , ALUopE , MemwriteE , ALUSrcE , RegwriteE , sign_extE;
    wire[25:0] target_E;
    wire[31:0] ALU_resultM , write_data;
    wire[1:0] rs_source , rt_source;
    wire[31:0] ALU_result;
    wire[2:0] Flag;
    wire[4:0] write_register;
    wire[4:0] write_registerM , write_registerW;
    wire MemreadM , MemtoRegM , MemwriteM , RegwriteM;
    wire[31:0] read_data_M2;
    wire[31:0] Memdata;
    wire MemtoRegW , RegwriteW;
    wire[31:0] ALU_resultW , MemdataW;
    reg CPU_enable;

    initial begin
        CPU_enable = 1;
    end

    PC_checker pc_checker(CLK , NEW_PC , BRC_PC , PC_BRCH_INTO , JUMP_TO_PC , JUMPSIGN , PC_write , PC);
    instruction_memory Instruction_memory(CLK , PC , ENABLE , NEW_PC , INSTRUCTION);
    enable_checker Enable_checker(INSTRUCTION , ENABLE);
    IF_ID_buffer IF_ID_Buffer(INSTRUCTION , NEW_PC , IF_flush , IF_ID_write , CLK , ENABLE , next_PC , instruction_F);
    decode Decode(instruction_F , opcode , rs , rt , rd , imme , funct , shamt , target);
    control_signal control_signal(opcode , funct , ID_EX_flush , zero_flag , RegDst , Branch , Memread , MemtoReg , ALUop , Memwrite , ALUSrc ,  Regwrite , sign_ext , IF_flush , PC_BRCH_INTO , JUMPSIGN);
    Register register_part(CLK , next_PC , write_back_data , write_registerW , RegwriteW , opcode , rs , rt , imme , target , read_data1 , read_data2 , BRC_PC , JUMP_TO_PC , zero_flag);
    hazard_unit Hazard_unit(rs , rt , rt_E , MemreadE , MemwriteE , PC_write , IF_ID_write , ID_EX_flush);
    ID_EX_buffer ID_EX_Buffer(
    CLK , read_data1 , read_data2 , rs , rt , rd , imme , opcode , shamt , funct , target , next_PC , 
    RegDst , Memread , MemtoReg , ALUop , Memwrite , ALUSrc , Regwrite , sign_ext ,
    RegDstE , MemreadE , MemtoRegE , ALUopE , MemwriteE , ALUSrcE , RegwriteE , sign_extE,
    read_data_E1 , read_data_E2 , imme_E , rs_E , rt_E , rd_E , opcode_E , shamt_E , funct_E , target_E , next_PC_E);
    ALU  ALU_part(
    opcode_E , shamt_E , funct_E , next_PC_E ,  read_data_E1 , read_data_E2 , ALU_resultM , write_back_data , imme_E , sign_extE, rs_source , rt_source , ALUSrcE , Flag , ALU_result );
    Write_register_checker Write_register(opcode_E , rt_E , rd_E , RegDstE , write_register);
    forwarding_unit Forwarding(CLK , rs_E , rt_E , write_registerM , write_registerW , RegwriteM , RegwriteW , rs_source , rt_source);
    EX_MEM_buffer EX_MEM_Buffer(CLK , ALU_result , MemreadE , MemtoRegE , MemwriteE , RegwriteE , write_register , read_data_E2 , 
                                      ALU_resultM , MemreadM , MemtoRegM , MemwriteM , RegwriteM , write_registerM , read_data_M2);
    MainMemory MainMEMORY(ALU_resultM , read_data_M2 , MemreadM , MemwriteM , Memdata);
    MEM_WB_buffer MEM_WB_Buffer(CLK , MemtoRegM , RegwriteM , write_registerM , ALU_resultM , Memdata,
                                      MemtoRegW , RegwriteW , write_registerW , ALU_resultW , MemdataW);
    Check_write_back_data check_write_back_data(MemtoRegW , ALU_resultW , MemdataW , write_back_data);

    integer i;
    integer j;
    integer k;
    integer fp_w;
    // initial begin
    //     $dumpfile("test.vcd");
    //     $dumpvars(0 , pc , pc_checker , Instruction_memory , Enable_checker , IF_ID_Buffer , Decode , control_signal , register_part , ID_EX_Buffer ,  ALU_part , Write_register , EX_MEM_Buffer , MainMEMORY , MEM_WB_Buffer , check_write_back_data , Forwarding , Hazard_unit);
    // end
    always @(INSTRUCTION) begin
        if(INSTRUCTION == 32'b11111111111111111111111111111111) begin
            CPU_enable <= 0;
        end
    end
    always @(CPU_enable) begin
        if(CPU_enable == 0) begin
            fp_w=$fopen("data.bin","w");
            #40;
            for (j=0; j < 512; j = j + 1) begin
                $display("%b", MainMEMORY.DATA_RAM[j]);
                $fwrite(fp_w, "%b\n",MainMEMORY.DATA_RAM[j]);
            end
            $finish();
        end
    end
endmodule
